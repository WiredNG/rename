package WiredRenameBitmap;

import GetPut::*;
import FIFOF::*;
import PriorityEncodeOH::*;

interface WiredRenameBitmap;
endinterface

module mkWiredRenameBitmap(

);

endmodule

endpackage